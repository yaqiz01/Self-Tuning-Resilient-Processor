LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY razor_latch IS
PORT ( input : IN STD_LOGIC_VECTOR(31 downto 0);
   write_enable :IN STD_LOGIC;
   clock: IN STD_LOGIC;
   reset: IN STD_LOGIC;
   output : OUT STD_LOGIC_VECTOR(31 downto 0);
   shadow_out: OUT STD_LOGIC_VECTOR(31 downto 0);
   restore: out std_logic );
END razor_latch;

ARCHITECTURE structure OF razor_latch IS

component reg_32
PORT ( input : IN STD_LOGIC_VECTOR(31 downto 0);
   write_enable :IN STD_LOGIC;
   clock: IN STD_LOGIC;
   reset: IN STD_LOGIC;
   output : OUT STD_LOGIC_VECTOR(31 downto 0)
   );
END component;

component comparator_32
PORT ( data_operandA, data_operandB     : IN STD_LOGIC_VECTOR(31 downto 0);
	not_equal: out std_logic;
	less_than: out std_logic);
END component;

component razor_dflipflop
   port
   ( clock, reset,data,restore_data : in std_logic;
   enable : in  STD_LOGIC_VECTOR(1 downto 0);
      output : out std_logic;
      restore: out std_logic
   );
end component;

signal main_ff_out: STD_LOGIC_VECTOR(31 downto 0);
signal shadow_latch_out: STD_LOGIC_VECTOR(31 downto 0);
signal enable_comb: STD_LOGIC_VECTOR(1 downto 0);
signal main_shadow_equal: std_logic;
signal noteq_rising_edge: std_logic;

BEGIN
enable_comb(0) <= main_shadow_equal when noteq_rising_edge = '0' else '0';
enable_comb(1) <= write_enable;

d0: razor_dflipflop port map(clock,reset,input(0),shadow_latch_out(0),enable_comb,main_ff_out(0),noteq_rising_edge);

G1: for i in 31 downto 1 generate
	d31_1: razor_dflipflop port map(clock,reset,input(i),shadow_latch_out(i),enable_comb,main_ff_out(i),open);
end generate;

shadow_latch: reg_32 port map (input, write_enable, not clock, reset, shadow_latch_out);
comparator: comparator_32 port map(main_ff_out,shadow_latch_out,main_shadow_equal,open);
output <= main_ff_out;
shadow_out <= shadow_latch_out;
restore <= noteq_rising_edge;

END structure;
